`include "def.v"

/*
    指令只读存储器ROM
*/
module InstMem(
    input wire ce, //读使能信号，来自IF的romCe
    input wire[31:0] addr, //读地址信号，来自IF的PC
    output reg[31:0] data //读取的指令，流入IF
);
    //1024个32位寄存器
    reg[31:0] ROM[1023:0]; 

    //组合逻辑语句块，按字读取指令
    always@(*)
    begin
        if(ce == `ROMCE_ENABLE)
            data <= ROM[addr[11:2]];
        else
            data <= 32'b0;
    end

    //ROM中预先存储的指令字
    initial
    begin
/*      
        //initial
        ROM[0] <= 32'h3463000a;
        ROM[1] <= 32'h34840001;
        ROM[2] <= 32'h34210000;
        ROM[3] <= 32'h0c000006;
        ROM[4] <= 32'h8c060004;
        ROM[5] <= 32'h00000000;
        ROM[6] <= 32'h00441020;
        ROM[7] <= 32'h20840001;
        ROM[8] <= 32'hac220000;
        ROM[9] <= 32'h20210004;
        ROM[10] <= 32'h1483fffb;
        ROM[11] <= 32'h03e00008;
*/


        //mul-div
        ROM[0] <= 32'h34011100; //ori r1, r0 0x1100 r1 = 00001100
        ROM[1] <= 32'h34020020; //ori r2, r0 0x0020 r2 = 00000020
        ROM[2] <= 32'b00000_00010_00000_00000_00000_011001; //multu r1,r2  22000
        ROM[3] <= 32'h3403ffff; //roi r3, r0, 0xffff r3 = 0000ffff
        ROM[4] <= 32'b00000_00000_00011_00011_10000_000000; //sll  r3, r3, 0x10 r3 = ffff0000
        ROM[5] <= 32'b00000_00011_00010_00000_00000_011000; //mult r3, r2  lo = ffe00000 hi = ffffffff
        ROM[6] <= 32'b00000_00001_00010_00000_00000_011011; //div  r1,r2   lo = 88h      hi = 0
        ROM[7] <= 32'b00000_00011_00010_00000_00000_011010; //divu r3, r2  lo = ffffff80 hi = 0


        //ori R0,1100 -- R1 --00001100
        //ROM[0] = 32'h34011100;
	//ori R0,0020 -- R2 --00000020
        //ROM[1] = 32'h34020020;
	//ori R0,ff00 -- R3 --0000ff00
        //ROM[2] = 32'h3403ff00;
	//ori R0,ffff -- R4 --0000ffff
        //ROM[3] = 32'h3404ffff;
		
	//I?????
/*
	//andi R0,ffff --R5 --00000000
	ROM[4] = 32'h3005ffff;
	//xori R0,ffff --R6 --0000ffff
	ROM[5] = 32'h3806ffff;
	//addi R0,ffff --R7 --ffffffff
	ROM[6] = 32'h2007ffff;
	//subi R0,ffff --R8 --00000001
	ROM[7] = 32'h2408ffff;
	//lui  R0,ffff --R9 --ffff0000
	ROM[8] = 32'h3C09ffff;
*/
		
	//R1=00001100 R2=00000020
	//ROM[4] = 32'b000000_00001_00010_00101_00000_100000;//add,R5,R1,R2  00001120
	//ROM[5] = 32'b000000_00001_00010_00110_00000_100101;//or,R6,R1,R2   00001120

	//R?????

	//ROM[6] = 32'b000000_00001_00010_00111_00000_100010;//sub,R7,R1,R2  000010e0
	//ROM[7] = 32'b000000_00001_00010_01000_00000_100100;//and,R8,R1,R2  00000000
	//ROM[8] = 32'b000000_00001_00010_01001_00000_100110;//xor,R9,R1,R2  00001120

	//lui  R0,ffff --R10 --ffff0000
	//ROM[9] = 32'h3C0Affff;

		
	//R11=fffe0000 R12=7fff8000  R13=ffff8000
	// Ra=sa={25'b0,imm[10:6]}
	//ROM[10] = 32'b000000_00000_01010_01011_00001_000000;//sll,R11,Ra,R10
	//ROM[11] = 32'b000000_00000_01010_01100_00001_000010;//srl,R12,Ra,R10  		
	//ROM[12] = 32'b000000_00000_01010_01101_00001_000011;//sra,R13,Ra,R10
        //ROM[6] = 32'b000000_00010_00001_00111_00000_101010;//slt,R7<-(R2<R1),signed

	//J- JR?????

	//ROM[6] = 32'h18000000;  //j 0		??000110
	//ROM[6] = 32'h14000000; //jal 0		??000101
	//ROM[6] = 32'h34070000;//ori,R7,0000
	//ROM[7] = 32'b000000_00111_00000_00000_001000; //jr R7		??001000 
	//ROM[7] = 32'b000000_00111_00000_00000_001001; //jalr R0		??001001


	//J+?????
	//R1=00001100 R2=00000020 R3=000000ff R4=0000ffff R5=00001120 R6=00001120
	//ROM[6] = 32'b010000_00101_00110_0000_0000_0000_0000;  //beq r5,r6,0 		??010000
	//ROM[6] = 32'b010001_00001_00110_0000_0000_0000_0000;  //bne r5,r6,0 		??010001
	//ROM[6] = 32'b000111_00010_00000_0000_0000_0000_0000;  //bltz r2,0 		??010010
	//ROM[6] = 32'b000001_00001_00000_0000_0000_0000_0000;  //bgtz r1,0 		??010011

        //mf/mthi,mf/mtlo
        ROM[8] = 32'h000000_00000_00000_01000_00000_010000;  //R8 <- hi
        ROM[9] = 32'h000000_00000_00000_01001_00000_010010;  //R9 <- lo
        ROM[10] = 32'h000000_01000_00000_00000_00000_010001; //hi <- R8
        ROM[11] = 32'h000000_01001_00000_00000_00000_010011; //lo <- R9

/*
        ROM[0] = 32'h3401ffff;
        ROM[1] = 32'h3402ffff;
        ROM[2] = 32'h3403ffff;
        ROM[3] = 32'h3404ffff;
        ROM[4] = 32'h0000000c;  //syscall??
        ROM[5] = 32'h3405ffff;
        ROM[6] = 32'h3406ffff;
        ROM[16] = 32'h340affff;  //??????????
        ROM[17] = 32'h340bffff;
        ROM[18] = 32'h42000018;  //eret??
        //???????????mtc????Status????IM???IE??
        //???????????????
        ROM[0] = 32'h34020000;   //ori $2, $0, 0
        ROM[1] = 32'h34010014;   //ori $1, $0, 20
        ROM[2] = 32'h40815800;   //mtc0 $1, $11 set compare=20
        ROM[3] = 32'h3c011000;   //lui $1, 0x1000
        ROM[4] = 32'h34210401;   //ori $1, $1, 0x0401
        ROM[5] = 32'h40816000;   //mtc0 $1, $12 set status,enable int
        ROM[6] =32'h08000006;   //lpt: j lpt
        //interproc first addr 0x0050
        ROM[20] = 32'h34030001;   //ORI $3, $0, 1
        ROM[21] = 32'h34040014;   //ORI $4, $0, 20
        ROM[22] = 32'h00431020;   //ADD $2, $2, $3
        ROM[23] = 32'h40015800;   //MFC $1, $11  read compare
        ROM[24] = 32'h00240820;   //ADD $1, $1, $4
        ROM[25] = 32'h40815800;   //MTC0 $1, $11 set compare
        ROM[26] = 32'h42000018;   //eret
*/

    end
endmodule

//独立测试模块
module InstMem_tb;
    reg ce;
    reg[31:0] addr;
    wire[31:0] data;

    InstMem U1(ce,addr,data);

    initial
    begin
        addr <= 32'b0;
        ce <= `RST_ENABLE;

    #10 ce <= `RST_DISABLE;
    #5  $stop;
    end

    always #1 addr <= addr + 4;

endmodule